DataMemory.v                                                                                        0000644 0001750 0001750 00000005153 14763111070 011405  0                                                                                                    ustar   ben                             ben                                                                                                                                                                                                                    `timescale 1ns / 1ps

`define SIZE 1024

module DataMemory(ReadData , Address , WriteData , MemoryRead , MemoryWrite , Clock);
   input [63:0]      WriteData;
   input [63:0]      Address;
   input             Clock, MemoryRead, MemoryWrite;
   output reg [63:0] ReadData;

   reg [7:0] 	     memBank [`SIZE-1:0];


   // This task is used to write arbitrary data to the Data Memory by
   // the intialization block.
   task initset;
      input [63:0] addr;
      input [63:0] data;
      begin
	 memBank[addr] =  data[63:56] ; // Big-endian for the win...
	 memBank[addr+1] =  data[55:48];
	 memBank[addr+2] =  data[47:40];
	 memBank[addr+3] =  data[39:32];
	 memBank[addr+4] =  data[31:24];
	 memBank[addr+5] =  data[23:16];
	 memBank[addr+6] =  data[15:8];
	 memBank[addr+7] =  data[7:0];
      end
   endtask


   initial
     begin
        // preseting some data in the data memory used by test #1

        // Address 0x0 gets 0x1
        initset( 64'h0,  64'h1);  //Counter variable
        initset( 64'h8,  64'ha);  //Part of mask
        initset( 64'h10, 64'h5);  //Other part of mask
        initset( 64'h18, 64'h0ffbea7deadbeeff); //big constant
        initset( 64'h20, 64'h0); //clearing space

        // Add any data you need for your tests here.

     end

   // This always block reads the data memory and places a double word
   // on the ReadData bus.
   always @(posedge Clock)
     begin
        if(MemoryRead)
          begin
             ReadData[63:56] <=  memBank[Address];
             ReadData[55:48] <=  memBank[Address+1];
             ReadData[47:40] <=  memBank[Address+2];
             ReadData[39:32] <=  memBank[Address+3];
             ReadData[31:24] <=  memBank[Address+4];
             ReadData[23:16] <=  memBank[Address+5];
             ReadData[15:8] <=  memBank[Address+6];
             ReadData[7:0] <=  memBank[Address+7];
          end
     end

   // This always block takes data from the WriteData bus and writes
   // it into the DataMemory.
   always @(posedge Clock)
     begin
        if(MemoryWrite)
          begin
             memBank[Address] <= #3 WriteData[63:56] ;
             memBank[Address+1] <= #3 WriteData[55:48];
             memBank[Address+2] <= #3 WriteData[47:40];
             memBank[Address+3] <= #3 WriteData[39:32];
             memBank[Address+4] <= #3 WriteData[31:24];
             memBank[Address+5] <= #3 WriteData[23:16];
             memBank[Address+6] <= #3 WriteData[15:8];
             memBank[Address+7] <= #3 WriteData[7:0];
             // Could be useful for debugging:
             // $display("Writing Address:%h Data:%h",Address, WriteData);
          end
     end
endmodule
                                                                                                                                                                                                                                                                                                                                                                                                                     InstructionMemory.v                                                                                 0000644 0001750 0001750 00000003546 14763111070 013061  0                                                                                                    ustar   ben                             ben                                                                                                                                                                                                                    `timescale 1ns / 1ps
/*
 * Module: InstructionMemory
 *
 * Implements read-only instruction memory
 * 
 */
module InstructionMemory(Data, Address);
   parameter T_rd = 20;
   parameter MemSize = 40;
   
   output [31:0] Data;
   input [63:0]  Address;
   reg [31:0] 	 Data;
   
   /*
    * ECEN 350 Processor Test Functions
    * Texas A&M University
    */
   
   always @ (Address) begin

      case(Address)

	/* Test Program 1:
	 * Program loads constants from the data memory. Uses these constants to test
	 * the following instructions: LDUR, ORR, AND, CBZ, ADD, SUB, STUR and B.
	 * 
	 * Assembly code for test:
	 * 
	 * 0: LDUR X9, [XZR, 0x0]    //Load 1 into x9
	 * 4: LDUR X10, [XZR, 0x8]   //Load a into x10
	 * 8: LDUR X11, [XZR, 0x10]  //Load 5 into x11
	 * C: LDUR X12, [XZR, 0x18]  //Load big constant into x12
	 * 10: LDUR X13, [XZR, 0x20]  //load a 0 into X13
	 * 
	 * 14: ORR X10, X10, X11  //Create mask of 0xf
	 * 18: AND X12, X12, X10  //Mask off low order bits of big constant
	 * 
	 * loop:
	 * 1C: CBZ X12, end  //while X12 is not 0
	 * 20: ADD X13, X13, X9  //Increment counter in X13
	 * 24: SUB X12, X12, X9  //Decrement remainder of big constant in X12
	 * 28: B loop  //Repeat till X12 is 0
	 * 2C: STUR X13, [XZR, 0x20]  //store back the counter value into the memory location 0x20
	 */
	

	63'h000: Data = 32'hF84003E9;
	63'h004: Data = 32'hF84083EA;
	63'h008: Data = 32'hF84103EB;
	63'h00c: Data = 32'hF84183EC;
	63'h010: Data = 32'hF84203ED;
	63'h014: Data = 32'hAA0B014A;
	63'h018: Data = 32'h8A0A018C;
	63'h01c: Data = 32'hB400008C;
	63'h020: Data = 32'h8B0901AD;
	63'h024: Data = 32'hCB09018C;
	63'h028: Data = 32'h17FFFFFD;
	63'h02c: Data = 32'hF80203ED;
	63'h030: Data = 32'hF84203ED;  //One last load to place stored value on memdbus for test checking.

	/* Add code for your tests here */

	
	default: Data = 32'hXXXXXXXX;
      endcase
   end
endmodule
                                                                                                                                                          Mux21.v                                                                                             0000644 0001750 0001750 00000000603 14773762004 010264  0                                                                                                    ustar   ben                             ben                                                                                                                                                                                                                    module Mux21(out, in,  sel);
   // declare ports & internal wires
   input [1:0] in;
   input       sel;
   output      out;
   wire	       w1, w2, w3;

   // instantiate logic gates
   not not1(w1, sel); // w1 = sel'
   and and1(w2, in[0], w1); // w2 = (in[0])*sel'
   and and2(w3, in[1], sel); // w3 = (in[1])*sel
   or or1(out, w2, w3); // out = (in[1]*sel) + (in[0]*sel')

endmodule
                                                                                                                             NextPClogic.v                                                                                       0000644 0001750 0001750 00000001152 14771527055 011532  0                                                                                                    ustar   ben                             ben                                                                                                                                                                                                                    module NextPClogic(NextPC, CurrentPC, SignExtImm64, Branch, ALUZero, Uncondbranch); 
   input [63:0] CurrentPC, SignExtImm64; 
   input 	Branch, ALUZero, Uncondbranch; 
   output reg [63:0] NextPC; 

   always @(*)
     begin
	// Check branch conditions; if branch not taken, PC += 4
	     if (Uncondbranch) // unconditional branch taken
	       NextPC = CurrentPC + (SignExtImm64 << 2);
	     else  if (Branch && ALUZero) // conditional branch taken
	       NextPC = CurrentPC + (SignExtImm64 << 2);
	     else // neither path taken, PC += 4
	       NextPC = CurrentPC + 64'b100;
     end // always @ (*)


endmodule
                                                                                                                                                                                                                                                                                                                                                                                                                      RegisterFile.v                                                                                      0000644 0001750 0001750 00000001662 14771535110 011734  0                                                                                                    ustar   ben                             ben                                                                                                                                                                                                                    `timescale 1ns/1ps
module RegisterFile(BusA, BusB, BusW, RA, RB, RW, RegWr, Clk);
output [63:0] BusA; //64 bit wide buses
output [63:0] BusB;
input [63:0] BusW;
input [4:0] RA; //5-bit wide register indexes
input [4:0] RB;
input [4:0] RW;
input RegWr; //write enable
input Clk;


reg [63:0] registers [31:0]; //internal register file

//initial begin
//   registers[31] = 64'b0; //set register 31 to be 0
//end

assign #2  BusA = (RA == 5'b11111) ? 64'b0 : registers[RA]; //assigning BusA with contents in RegisterA after 2 sec delay
assign #2  BusB = (RB == 5'b11111) ? 64'b0 : registers[RB]; //assigning BusB with contents in RegisterB after 2 sec delay


always@(negedge Clk) begin //writing to a register on falling clock edge
	if (RegWr && !(RW == 5'b11111)) //checking if Write is enabled (do not allow writing to register 31)
	  registers[RW] <= #3 BusW; //writing BusW contents to register
	
end


endmodule
                                                                              SignExtender.v                                                                                      0000644 0001750 0001750 00000001760 14767303403 011751  0                                                                                                    ustar   ben                             ben                                                                                                                                                                                                                    module SignExtender(BusImm, Inst, Ctrl);
   // declare i/o ports 
   output reg [63:0] BusImm; 
   input [25:0]  Inst; 
   input [1:0]	 Ctrl;

   // For I-type: Ctrl = [0, 0]
   // For D-type: Ctrl = [0, 1]
   // For B-type: Ctrl = [1, 0]
   // For CB-type: Ctrl = [1, 1]

   // switch over all possibilities of Ctrl
    always @(*)
      begin

       case (Ctrl)
         2'b00:  BusImm = {{52{1'b0}}, Inst[21:10]}; //zero extending 12 bit immediate stored in I[21:10] since this is R-type
         2'b01:  BusImm = {{55{Inst[20]}}, Inst[20:12]}; //sign extending 9 bit immediate stored in I[20:12] since this is D-type (memory access)
         2'b10:  BusImm = {{38{Inst[25]}}, Inst[25:0]}; //sign extending 26 bit immediate stored in I[25:0] since this is B-type (unconditional branch)
         2'b11:  BusImm = {{52{Inst[23]}}, Inst[23:5]}; //sign extending 19 bit immediate stored in I[23:5] since this is CB-type (conditional branch)
	 default: BusImm = 0;
       endcase

      end
   
   
endmodule
                SingleCycleControl.v                                                                                0000644 0001750 0001750 00000013514 14773767353 013133  0                                                                                                    ustar   ben                             ben                                                                                                                                                                                                                    `define OPCODE_ANDREG 11'b?0001010???
`define OPCODE_ORRREG 11'b?0101010???
`define OPCODE_ADDREG 11'b?0?01011???
`define OPCODE_SUBREG 11'b?1?01011???

`define OPCODE_ADDIMM 11'b?0?10001???
`define OPCODE_SUBIMM 11'b?1?10001???

`define OPCODE_MOVZ   11'b110100101??

`define OPCODE_B      11'b?00101?????
`define OPCODE_CBZ    11'b?011010????

`define OPCODE_LDUR   11'b??111000010
`define OPCODE_STUR   11'b??111000000

module control(
	       output reg 	reg2loc,
	       output reg 	alusrc,
	       output reg 	mem2reg,
	       output reg 	regwrite,
	       output reg 	memread,
	       output reg 	memwrite,
	       output reg 	branch,
	       output reg 	uncond_branch,
	       output reg [3:0] aluop,
	       output reg [1:0] signop,
	       input [10:0] 	opcode
	       );

   always @(*)
     begin
	casez (opcode)

          /* Add cases here for each instruction your processor supports */
	  `OPCODE_ANDREG: // AND operation (R-type)
	    begin
               reg2loc       = 1'b0;
               alusrc        = 1'b0;
               mem2reg       = 1'b0;
               regwrite      = 1'b1;
               memread       = 1'b0;
               memwrite      = 1'b0;
               branch        = 1'b0;
               uncond_branch = 1'b0;
               aluop         = 4'b0000;
               signop        = 2'bxx;
            end // case: `OPCODE_ANDREG

	  `OPCODE_ORRREG: // OR (R-type)
	    begin
               reg2loc       = 1'b0;
               alusrc        = 1'b0;
               mem2reg       = 1'b0;
               regwrite      = 1'b1;
               memread       = 1'b0;
               memwrite      = 1'b0;
               branch        = 1'b0;
               uncond_branch = 1'b0;
               aluop         = 4'b0001;
               signop        = 2'bxx;
            end // case: `OPCODE_ORREG

	    `OPCODE_ADDREG: // ADD (R-type)
	    begin
               reg2loc       = 1'b0;
               alusrc        = 1'b0;
               mem2reg       = 1'b0;
               regwrite      = 1'b1;
               memread       = 1'b0;
               memwrite      = 1'b0;
               branch        = 1'b0;
               uncond_branch = 1'b0;
               aluop         = 4'b0010;
               signop        = 2'bxx;
            end // case: `OPCODE_ADDREG

	    `OPCODE_SUBREG: // SUB (R-type)
	    begin
               reg2loc       = 1'b0;
               alusrc        = 1'b0;
               mem2reg       = 1'b0;
               regwrite      = 1'b1;
               memread       = 1'b0;
               memwrite      = 1'b0;
               branch        = 1'b0;
               uncond_branch = 1'b0;
               aluop         = 4'b0110;
               signop        = 2'bxx;
            end // case: `OPCODE_SUBREG

	    `OPCODE_ADDIMM: // ADD (I-type)
	    begin
               reg2loc       = 1'bx;
               alusrc        = 1'b1;
               mem2reg       = 1'b0;
               regwrite      = 1'b1;
               memread       = 1'b0;
               memwrite      = 1'b0;
               branch        = 1'b0;
               uncond_branch = 1'b0;
               aluop         = 4'b0010;
               signop        = 2'b00;
            end // case: `OPCODE_ADDIMM

	  `OPCODE_SUBIMM: // SUB (I-type)
	    begin
               reg2loc       = 1'bx;
               alusrc        = 1'b1;
               mem2reg       = 1'b0;
               regwrite      = 1'b1;
               memread       = 1'b0;
               memwrite      = 1'b0;
               branch        = 1'b0;
               uncond_branch = 1'b0;
               aluop         = 4'b0110;
               signop        = 2'b00;
	    end // case: `OPCODE_SUBIMM

	 `OPCODE_B: // Branch (B-type)
	    begin
               reg2loc       = 1'bx;
               alusrc        = 1'bx;
               mem2reg       = 1'b0;
               regwrite      = 1'b0;
               memread       = 1'b0;
               memwrite      = 1'b0;
               branch        = 1'bx;
               uncond_branch = 1'b1;
               aluop         = 4'bxxxx;
               signop        = 2'b10;
	    end // case: `OPCODE_B

	  `OPCODE_CBZ: // CBZ (CB-type)
	    begin
               reg2loc       = 1'b1;
               alusrc        = 1'b0;
               mem2reg       = 1'b0;
               regwrite      = 1'b0;
               memread       = 1'b0;
               memwrite      = 1'b0;
               branch        = 1'b1;
               uncond_branch = 1'b0;
               aluop         = 4'b0111;
               signop        = 2'b11;
	    end // case: `OPCODE_CBZ

	  `OPCODE_LDUR: // LDUR (D-type)
	    begin
               reg2loc       = 1'bx;
               alusrc        = 1'b1;
               mem2reg       = 1'b1;
               regwrite      = 1'b1;
               memread       = 1'b1;
               memwrite      = 1'b0;
               branch        = 1'b0;
               uncond_branch = 1'b0;
               aluop         = 4'b0010;
               signop        = 2'b01;
	    end // case: `OPCODE_LDUR

	  `OPCODE_STUR: // STUR (D-type)
	    begin
               reg2loc       = 1'b1;
               alusrc        = 1'b1;
               mem2reg       = 1'b0;
               regwrite      = 1'b0;
               memread       = 1'b0;
               memwrite      = 1'b1;
               branch        = 1'b0;
               uncond_branch = 1'b0;
               aluop         = 4'b0010;
               signop        = 2'b01;
	    end // case: `OPCODE_STUR

	  /* Add support for MOVZ */
	  

          default:
            begin
               reg2loc       = 1'bx;
               alusrc        = 1'bx;
               mem2reg       = 1'bx;
               regwrite      = 1'b0;
               memread       = 1'b0;
               memwrite      = 1'b0;
               branch        = 1'b0;
               uncond_branch = 1'b0;
               aluop         = 4'bxxxx;
               signop        = 2'bxx;
            end
	endcase
     end

endmodule

                                                                                                                                                                                    SingleCycleProcTest.v                                                                               0000644 0001750 0001750 00000006027 14773766131 013250  0                                                                                                    ustar   ben                             ben                                                                                                                                                                                                                    `timescale 1ns / 1ps

`define STRLEN 32
`define HalfClockPeriod 60
`define ClockPeriod `HalfClockPeriod * 2

module SingleCycleProcTest_v;

   initial
     begin
        $dumpfile("singlecycle.vcd");
        $dumpvars;
     end

   // These tasks are used to check if a given test has passed and
   // confirm that all tests passed.
   task passTest;
      input [63:0] actualOut, expectedOut;
      input [`STRLEN*8:0] testType;
      inout [7:0] 	  passed;

      if(actualOut == expectedOut) begin $display ("%s passed", testType); passed = passed + 1; end
      else $display ("%s failed: 0x%x should be 0x%x", testType, actualOut, expectedOut);
   endtask

   task allPassed;
      input [7:0] passed;
      input [7:0] numTests;

      if(passed == numTests) $display ("All tests passed");
      else $display("Some tests failed: %d of %d passed", passed, numTests);
   endtask

   // Inputs
   reg 		  CLK;
   reg 		  Reset_L;
   reg [63:0] 	  startPC;
   reg [7:0] 	  passed;
   reg [15:0] 	  watchdog;

   // Outputs
   wire [63:0] 	  MemtoRegOut;
   wire [63:0] 	  currentPC;

   // Instantiate the Unit Under Test (UUT)
   singlecycle uut (
		    .CLK(CLK),
		    .resetl(Reset_L),
		    .startpc(startPC),
		    .currentpc(currentPC),
		    .MemtoRegOut(MemtoRegOut)
		    );

   initial begin
      // Initialize Inputs
      Reset_L = 1;
      startPC = 0;
      passed = 0;

      // Initialize Watchdog timer
      watchdog = 0;

      // Wait for global reset
      #(1 * `ClockPeriod);

      // Program 1
      #1
        Reset_L = 0; startPC = 0;
      @(posedge CLK);
      @(negedge CLK);
      @(posedge CLK);
      Reset_L = 1;

      // ***********************************************************
      // This while loop will continue cycling the processor until the
      // PC reaches the final instruction in the first test.  If the
      // program forms an infinite loop, never reaching the end, the
      // watchdog timer will kick in and kill simulation after 64K
      // cycles.
      // ***********************************************************

      while (currentPC < 64'h30)
        begin
	   @(posedge CLK);
	   @(negedge CLK);
           $display("CurrentPC:%h",currentPC);
        end
      passTest(MemtoRegOut, 64'hF, "Results of Program 1", passed);

      // ***********************************************************
      // Add your new tests here
      // ***********************************************************

      // Done
      allPassed(passed, 1);   // Be sure to change the one to match
      // the number of tests you add.
      $finish;
   end

   // Initialize the clock to be 0
   initial begin
      CLK = 0;
   end

   // The following is correct if clock starts at LOW level at StartTime //
   always begin
      #`HalfClockPeriod CLK = ~CLK;
      #`HalfClockPeriod CLK = ~CLK;
      watchdog = watchdog +1;
   end

   // Kill the simulation if the watchdog hits 64K cycles
   always @*
     if (watchdog == 16'hFF)
       begin
          $display("Watchdog Timer Expired.");
          $finish;
       end


endmodule

                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         SingleCycleProc.v                                                                                   0000644 0001750 0001750 00000007001 14773765455 012411  0                                                                                                    ustar   ben                             ben                                                                                                                                                                                                                    module singlecycle(
		   input 	     resetl,
		   input [63:0]      startpc,
		   output reg [63:0] currentpc,
		   output [63:0]     MemtoRegOut,  // this should be
						   // attached to the
						   // output of the
						   // MemtoReg Mux
		   input 	     CLK
		   );

   // Next PC connections
   wire [63:0] 			     nextpc;       // The next PC, to be updated on clock cycle

   // Instruction Memory connections
   wire [31:0] 			     instruction;  // The current instruction

   // Parts of instruction
   wire [4:0] 			     rd;            // The destination register
   wire [4:0] 			     rm;            // Operand 1
   wire [4:0] 			     rn;            // Operand 2
   wire [10:0] 			     opcode;

   // Control wires
   wire 			     reg2loc;
   wire 			     alusrc;
   wire 			     mem2reg;
   wire 			     regwrite;
   wire 			     memread;
   wire 			     memwrite;
   wire 			     branch;
   wire 			     uncond_branch;
   wire [3:0] 			     aluctrl;
   wire [1:0] 			     signop;

   // Register file connections
   wire [63:0] 			     regoutA;     // Output A
   wire [63:0] 			     regoutB;     // Output B

   // ALU connections
   wire [63:0] 			     aluout;
   wire 			     zero;

   /* Add Multiplexer signal controlled by AluSrc */
   wire [63:0]			     alu_arg2;
   

   // Sign Extender connections
   wire [63:0]			     extimm;

   // Data memory connections
   wire [63:0]			     readdata;
   

   // PC update logic
   always @(negedge CLK)
     begin
        if (resetl)
          currentpc <= #3 nextpc;
        else
          currentpc <= #3 startpc;
     end

   // Parts of instruction
   assign rd = instruction[4:0];
   assign rm = instruction[9:5];
   assign rn = reg2loc ? instruction[4:0] : instruction[20:16];
   assign opcode = instruction[31:21];

   InstructionMemory imem(
			  .Data(instruction),
			  .Address(currentpc)
			  );

   control control(
		   .reg2loc(reg2loc),
		   .alusrc(alusrc),
		   .mem2reg(mem2reg),
		   .regwrite(regwrite),
		   .memread(memread),
		   .memwrite(memwrite),
		   .branch(branch),
		   .uncond_branch(uncond_branch),
		   .aluop(aluctrl),
		   .signop(signop),
		   .opcode(opcode)
		   );

   /*
    * Connect the remaining datapath elements below.
    * Do not forget any additional multiplexers that may be required.
    */

   // Instantiate data memory & connect ports
   DataMemory DataMem(
		      .ReadData(readdata),
		      .Address(aluout),
		      .WriteData(regoutB),
		      .MemoryRead(memread),
		      .MemoryWrite(memwrite),
		      .Clock(CLK)
		      );

   // Instantiate ALU & connect ports
   ALU Alu(
	   .BusW(aluout),
	   .BusA(regoutA),
	   .BusB(alu_arg2),
	   .ALUCtrl(aluctrl),
	   .Zero(zero)
	   );
   

   // Instantiate register file & connect ports
   RegisterFile RegFile(
			     .BusA(regoutA),
			     .BusB(regoutB),
			     .BusW(MemtoRegOut),
			     .RA(rm),
			     .RB(rn),
			     .RW(rd),
			     .RegWr(regwrite),
			     .Clk(CLK)
			     );

   // Instantiate sign extender & connect ports
   SignExtender SignExt(
			     .BusImm(extimm),
			     .Inst(instruction[25:0]),
			     .Ctrl(signop)
			     );

   // Instantiate the next PC logic
   NextPClogic PClogic(
			   .NextPC(nextpc),
			   .CurrentPC(currentpc),
			   .SignExtImm64(extimm),
			   .Branch(branch),
			   .ALUZero(zero),
			   .Uncondbranch(uncond_branch)
			   );


   // multiplex using control signal ALUSrc
   assign alu_arg2 = alusrc ? extimm : regoutB;

   // multiplex using control signal MemtoReg
   assign MemtoRegOut = mem2reg ? readdata : aluout;
   
   

endmodule

                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               